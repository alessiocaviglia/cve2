module vcve2_vrf_interface #(
    parameter int unsigned VLEN = 128,
    parameter int unsigned PIPE_WIDTH = 32
) (
    // Clock and Reset
    input   logic                       clk_i,
    input   logic                       rst_ni,

    // Read ports
    input   logic                       req_i,
    output  logic [PIPE_WIDTH-1:0]      rdata_a_o, rdata_b_o, rdata_c_o,

    // Write port
    input   logic [PIPE_WIDTH-1:0]      wdata_i,

    // Data memory interface
    output logic         data_req_o,
    input  logic         data_gnt_i,
    input  logic         data_rvalid_i,
    input  logic         data_err_i,
    input  logic         data_pmp_err_i,
    output logic         data_we_o,
    output logic [3:0]   data_be_o,
    output logic [31:0]  data_wdata_o,
    input  logic [31:0]  data_rdata_i,
    // LSU control signals
    output logic         data_load_addr_o,
    input  logic         lsu_gnt_i,

    // AGU
    output logic         agu_load_o,
    output logic         agu_get_rs1_o,
    output logic         agu_get_rs2_o,
    output logic         agu_get_rd_o,
    output logic         agu_incr_o,

    // ID signals
    input  logic [3:0]            sel_operation_i,    // each bit enables a different operation, 0 - R RS1, 1 - R RS2, 2 - R RS3, 3 - W RD
    input  logic                  memory_op_i,        // 0 - arithmetic operation, 1 - load/store operation
    input  logic                  interleaved_i,      // 0 - non-interleaved, 1 - interleaved
    output logic                  vector_done_o,      // signals the pipeline that the vector operation is finished (most likely with a write to the VRF)
    
    // LSU signals
    output logic                  lsu_req_o,          // signals the LSU that it can start the memory operation
    input  logic                  lsu_done_i,

    // CSR signals
    input vcve2_pkg::vlmul_e      lmul_i,
    input vcve2_pkg::vsew_e       sew_i,
    input logic [31:0]            vl_i
);

  import vcve2_pkg::*;

  parameter NUM_BYTE_OPS = (VLEN >> ($clog2(PIPE_WIDTH))) << 2; // (VLEN/PIPE_WIDTH) / 8 

  // VRF FSM signals
  vcve2_pkg::vrf_state_t vrf_state, vrf_next_state;
  logic [PIPE_WIDTH-3:0] num_iterations_q, num_iterations_d;
  logic [PIPE_WIDTH-1:0] num_bytes_elements;
  logic [1:0] offset_q, offset_d;
  logic first_iteration_d, first_iteration_q;
  logic last_iteration_d, last_iteration_q;
  logic [3:0] offset_be;
  logic no_offset;

  // Internal registers signals
  logic rs1_en, rs2_en, rs3_en, rd_en;    // rd is used only for load operations
  logic [PIPE_WIDTH-1:0] rs1_q, rs2_q, rs3_q, rd_q;
  logic [PIPE_WIDTH-1:0] rs1_d, rs2_d, rs3_d, rd_d;

  // Delayed grant for read operations in store
  logic read_delayed;
  logic curr_state_rdelay, next_state_rdelay;
  logic rdata_mux;
  logic rbuffer_en;
  logic [PIPE_WIDTH-1:0] rbuffer_q, rbuffer_d;
  // Delayed grant for write operations in interleaved
  logic write_delayed;
  logic curr_state_wdelay, next_state_wdelay;
  logic [1:0] wdata_mux;
  logic wbuffer_en, rd_buf_en;
  logic [PIPE_WIDTH-1:0] wbuffer_q, wbuffer_d;

  //////////////////
  // BE selector  //
  //////////////////

  // depending on vl we could need to access only a section of the 32 bit word
  always_comb begin
    no_offset = 1'b0;
    case (offset_q)
      2'b00: begin
        offset_be = 4'b0000;
        no_offset = 1'b1;
      end
      2'b01: offset_be = 4'b0001;
      2'b10: offset_be = 4'b0011;
      2'b11: offset_be = 4'b0111;
      default: offset_be = 4'b0000;
    endcase
  end
  // in interleaved operation the first read will not have the correct be but since it's only a read
  // it will not impact the state of the memory and the access will certainly be inside the vector register
  // since if there's an offset it means vl is certainly lower than vlmax
  assign data_be_o = (!no_offset && last_iteration_q) ? offset_be : 4'b1111;

  /////////////
  // VRF FSM //
  /////////////

  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      vrf_state <= VRF_IDLE;
      num_iterations_q <= '0;
      offset_q <= '0;
      first_iteration_q <= 1'b0;
      last_iteration_q <= 1'b0;
    end else begin
      vrf_state <= vrf_next_state;
      num_iterations_q <= num_iterations_d;
      offset_q <= offset_d;
      first_iteration_q <= first_iteration_d;
      last_iteration_q <= last_iteration_d;
    end
  end

  assign num_bytes_elements = vl_i<<sew_i;
  always_comb begin
    // register enables
    rs1_en = 1'b0;
    rs2_en = 1'b0;
    rs3_en = 1'b0;
    rd_en = 1'b0;
    write_delayed = 1'b0;
    read_delayed = 1'b0;
    // data memory interface
    data_req_o = 1'b0;
    data_we_o = 1'b0;
    // agu signals
    agu_load_o = 1'b0;
    agu_get_rs1_o = 1'b0;
    agu_get_rs2_o = 1'b0;
    agu_get_rd_o = 1'b0;
    agu_incr_o = 1'b0;
    // ID signals
    vector_done_o = 1'b0;
    num_iterations_d = num_iterations_q;
    offset_d = offset_q;
    first_iteration_d = first_iteration_q;
    last_iteration_d = last_iteration_q;
    // LSU signals
    lsu_req_o = 1'b0;
    data_load_addr_o = 1'b0;

    case (vrf_state)

      VRF_IDLE: begin
        last_iteration_d = 1'b0;
        // VRF stays idle until a request is made
        if (!req_i) begin
          vrf_next_state = VRF_IDLE;
          num_iterations_d = '0;
        // VRF receive a request
        end else begin
          // AGU - load addresses in the AGU
          agu_load_o = 1'b1;
          // Data memory if - load the start address
          if (memory_op_i) data_load_addr_o = 1'b1;
          // ITERATIONS COUNTER - we sample the correct value of num_iterations
          num_iterations_d = num_bytes_elements[31:2];
          offset_d = num_bytes_elements[1:0];
          vrf_next_state = VRF_START;
        end
      end

      VRF_START: begin
        // NEXT STATE SELECTION
        if (memory_op_i == 0) begin                   // ARITHMETIC OPERATION
          if (interleaved_i) begin                 // OPTIMIZED INTERLEAVED OPS
            first_iteration_d = 1'b1;
            data_req_o = 1'b1;                          // read RS1         
            agu_get_rs1_o = 1'b1;
            if (data_gnt_i) begin
              agu_incr_o = 1'b1;
              vrf_next_state = VRF_INT_READ1;
            end else vrf_next_state = VRF_START;
          end else begin                              // UNOPTIMIZED OPS
            if (sel_operation_i[0]) begin               // read RS1
              data_req_o = 1'b1;
              agu_get_rs1_o = 1'b1;
              if (data_gnt_i) begin
                agu_incr_o = 1'b1;
                vrf_next_state = VRF_READ1;
              end else vrf_next_state = VRF_START;
            end else if (sel_operation_i[1]) begin      // read RS2
              data_req_o = 1'b1;
              agu_get_rs2_o = 1'b1;
              if (data_gnt_i) begin
                agu_incr_o = 1'b1;
                vrf_next_state = VRF_READ2;
              end else vrf_next_state = VRF_START;
            end else if (sel_operation_i[3]) begin      // write RD
              data_we_o = 1'b1;
              data_req_o = 1'b1;
              agu_get_rd_o = 1'b1;
              if (data_gnt_i) begin
                agu_incr_o = 1'b1;
                vrf_next_state = VRF_WRITE;
              end else vrf_next_state = VRF_START;
            end else begin                              // illegal operation  
              vrf_next_state = VRF_IDLE;
            end
          end

        end else begin                                // MEMORY OPERATION
          first_iteration_d = 1'b1;
          if (sel_operation_i[2]==1'b1) begin           // store
            data_req_o = 1'b1;
            agu_get_rd_o = 1'b1;
            if (data_gnt_i) begin
              agu_incr_o = 1'b1;
              vrf_next_state = VRF_STORE_READ;
            end else vrf_next_state = VRF_START;
          end else if (sel_operation_i[3]==1'b1) begin  // load
            lsu_req_o = 1'b1;
            vrf_next_state = VRF_LOAD;
          end else begin                                // illegal operation
            vrf_next_state = VRF_IDLE;
          end
        end
        
      end

      /////////////////////////////////////////
      // Arithmetic operations - interleaved //
      /////////////////////////////////////////

      // In the following states the exit condition is the gnt signal since: gnt=1 => data_rvalid of the previous operation=1
      VRF_INT_READ1: begin
        // SAMPLE
        if (data_rvalid_i && !last_iteration_q) rs1_en = 1;
        // NEXT STATE SELECTION
        if (!first_iteration_q) begin
          data_we_o = 1'b1;
          data_req_o = 1'b1;
          agu_get_rd_o = 1'b1;
          if (data_gnt_i) begin
            write_delayed = 1'b0;
            agu_incr_o = 1'b1;
            vrf_next_state = VRF_INT_WRITE;
          end else begin
            write_delayed = 1'b1;
            vrf_next_state = VRF_INT_READ1;
          end
        end else begin
          first_iteration_d = 1'b0;
          vrf_next_state = VRF_INT_WRITE;
        end
      end

      VRF_INT_READ2: begin
        // SAMPLE
        if (data_rvalid_i) rs2_en = 1;
        // NEXT STATE SELECTION
        // if next operation is READ RD
        if (sel_operation_i[2]) begin
          data_req_o = 1'b1;
          agu_get_rd_o = 1'b1;
          if (data_gnt_i) begin
            vrf_next_state = VRF_INT_READ3;
          end else vrf_next_state = VRF_INT_READ2;
        // if next operation is WRITE RD
        end else if (sel_operation_i[3]) begin
          if (last_iteration_q) begin
            vrf_next_state = VRF_INT_READ1;
          end else begin
            data_req_o = 1'b1;
            agu_get_rs1_o = 1'b1;
            if (data_gnt_i) begin
              agu_incr_o = 1'b1;
              vrf_next_state = VRF_INT_READ1;
            end else vrf_next_state = VRF_INT_READ2;
          end
        // illegal operation
        end else begin
          vrf_next_state = VRF_IDLE;
        end
      end
      
      VRF_INT_READ3: begin
        // SAMPLE
        if (data_rvalid_i) rs3_en = 1;
        // NEXT STATE SELECTION
        if (sel_operation_i[3]) begin
          if (last_iteration_q) begin
            vrf_next_state = VRF_INT_READ1;
          end else begin
            data_req_o = 1'b1;
            agu_get_rs1_o = 1'b1;
            if (data_gnt_i) begin
              agu_incr_o = 1'b1;
              vrf_next_state = VRF_INT_READ1;
            end else vrf_next_state = VRF_INT_READ3;
          end
        // illegal operation
        end else begin
          vrf_next_state = VRF_IDLE;
        end
      end

      VRF_INT_WRITE: begin
        // NEXT STATE SELECTION - moving to the next iteration
        if (last_iteration_q) begin            // it's equal zero to take into account the first iteration
          vector_done_o = 1'b1;
          num_iterations_d = '0;
          vrf_next_state = VRF_IDLE;
        end else begin
          // if next operation is READ RS2
          if (sel_operation_i[1]) begin
            data_req_o = 1'b1;
            agu_get_rs2_o = 1'b1;
            if (data_gnt_i) begin
              agu_incr_o = 1'b1;
              if (num_iterations_q == (no_offset ? 1 : 0)) last_iteration_d = 1'b1;
              else num_iterations_d = num_iterations_q - 1;
              vrf_next_state = VRF_INT_READ2;
            end else begin
              num_iterations_d = num_iterations_q;   // if the operation wasn't accepted we need to repeat it
              vrf_next_state = VRF_INT_WRITE;
            end
          // illegal operation, go back to idle
          end else begin
            vrf_next_state = VRF_IDLE;
          end
        end
      end

      ///////////////////////////
      // Arithmetic operations //
      ///////////////////////////

      // In the following states the exit condition is the gnt signal since: gnt=1 => data_rvalid of the previous operation=1
      VRF_READ1: begin
        // SAMPLE
        if (data_rvalid_i) rs1_en = 1;
        // NEXT STATE SELECTION
        // from here we can only move to READ RS2
        if (sel_operation_i[1]) begin
          data_req_o = 1'b1;
          agu_get_rs2_o = 1'b1;
          if (data_gnt_i) begin
            agu_incr_o = 1'b1;
            vrf_next_state = VRF_READ2;
          end else vrf_next_state = VRF_READ1;
        end else begin
          vrf_next_state = VRF_IDLE;
        end
      end

      VRF_READ2: begin
        // SAMPLE
        if (data_rvalid_i) rs2_en = 1;
        // NEXT STATE SELECTION
        // if next operation is WRITE RD
        if (sel_operation_i[3]) begin
          data_we_o = 1'b1;
          data_req_o = 1'b1;
          agu_get_rd_o = 1'b1;
          if (data_gnt_i) begin
            agu_incr_o = 1'b1;
            vrf_next_state = VRF_WRITE;
          end else begin
            vrf_next_state = VRF_READ2;
          end
        end else begin
          // NEXT STATE SELECTION - moving to the next iteration
          if (num_iterations_q == 1) begin
            vector_done_o = 1'b1;
            num_iterations_d = '0;
            vrf_next_state = VRF_IDLE;
          end else begin
            num_iterations_d = num_iterations_q - 1;
            // if next operation is READ RS1
            if (sel_operation_i[0]) begin
              data_req_o = 1'b1;
              agu_get_rs1_o = 1'b1;
              if (data_gnt_i) begin
                agu_incr_o = 1'b1;
                vrf_next_state = VRF_READ1;
              end else begin
                num_iterations_d = num_iterations_q;   // if the operation wasn't accepted we need to repeat it
                vrf_next_state = VRF_READ2;
              end
            end else begin
              vrf_next_state = VRF_IDLE;
            end
          end
        end
      end

      VRF_WRITE: begin
        // NEXT STATE SELECTION - moving to the next iteration
        if (num_iterations_q == (no_offset ? 1 : 0)) begin
          vector_done_o = 1'b1;
          num_iterations_d = '0;
          vrf_next_state = VRF_IDLE;
        end else begin
          num_iterations_d = num_iterations_q - 1;
          // if next operation is READ RS2
          if (sel_operation_i[1]) begin
            data_req_o = 1'b1;
            agu_get_rs2_o = 1'b1;
            if (data_gnt_i) begin
              agu_incr_o = 1'b1;
              vrf_next_state = VRF_READ2;
            end else begin
              num_iterations_d = num_iterations_q;   // if the operation wasn't accepted we need to repeat it
              vrf_next_state = VRF_WRITE;
            end
          // if next operation is WRITE RD
          end else if (sel_operation_i[3]) begin
            data_we_o = 1'b1;
            data_req_o = 1'b1;
            agu_get_rd_o = 1'b1;
            if (data_gnt_i) begin
              agu_incr_o = 1'b1;
            end else begin
              num_iterations_d = num_iterations_q;   // if the operation wasn't accepted we need to repeat it
            end
            vrf_next_state = VRF_WRITE;
          end else begin
            vrf_next_state = VRF_IDLE;
          end
        end
      end

      ////////////////
      // Load/Store //
      ////////////////

      VRF_LOAD: begin
        if (lsu_done_i || last_iteration_q) begin
          // we sample only if it's not the last iteration
          if (lsu_done_i) rd_en = 1'b1;
          // we send a write request only if it's not the first iteration
          if (!first_iteration_q) begin
            data_we_o = 1'b1;
            data_req_o = 1'b1;
            agu_get_rd_o = 1'b1;
            if (data_gnt_i) begin
              agu_incr_o = 1'b1;
              vrf_next_state = VRF_LOAD_WRITE;
            end else begin
              write_delayed = 1'b1;
              vrf_next_state = VRF_LOAD_WAITGNT;
            end
          // if it's the first iteration we don't need to write the result
          end else begin
              first_iteration_d = 1'b0;
              vrf_next_state = VRF_LOAD_WRITE;
          end
        // we wait here for lsu to finish
        end else begin
          vrf_next_state = VRF_LOAD;
        end
      end

      // state where we wait for the grant from memory
      VRF_LOAD_WAITGNT: begin
        data_we_o = 1'b1;
        data_req_o = 1'b1;
        agu_get_rd_o = 1'b1;
        if (data_gnt_i) begin
          write_delayed = 1'b0;
          agu_incr_o = 1'b1;
          vrf_next_state = VRF_LOAD_WRITE;
        end else begin
          vrf_next_state = VRF_LOAD_WAITGNT;
        end
      end

      VRF_LOAD_WRITE: begin
        // if this is the last iteration we finish
        if (last_iteration_q) begin
          vector_done_o = 1'b1;
          num_iterations_d = '0;
          vrf_next_state = VRF_IDLE;
        // if the next iteration will be the last we don't need to read the operand
        end else if (num_iterations_q == (no_offset ? 1 : 0)) begin
          last_iteration_d = 1'b1;
          vrf_next_state = VRF_LOAD;
        // normal operation
        end else begin
          num_iterations_d = num_iterations_q - 1;
          lsu_req_o = 1'b1;
          vrf_next_state = VRF_LOAD;
        end
      end

      VRF_STORE_READ: begin
        // as soon as we see the value on the bus we sample it and tell the lsu it can proceed
        if (data_rvalid_i || last_iteration_q) begin
          if (data_rvalid_i) rs3_en = 1;
          if (!first_iteration_q) begin
            lsu_req_o = 1;
            if (!lsu_gnt_i) read_delayed = 1'b1;
          end
          vrf_next_state = VRF_STORE_WAITLSU;
        end else begin
          vrf_next_state = VRF_STORE_READ;
        end
      end

      VRF_STORE_WAITLSU: begin
        if (lsu_done_i || first_iteration_q) begin
          first_iteration_d = 1'b0;
          read_delayed = 1'b0;
          // Exit condition
          if (last_iteration_q) begin
            vector_done_o = 1'b1;
            num_iterations_d = '0;
            vrf_next_state = VRF_IDLE;
          // In the last cycle we don't read the operand
          end else if (num_iterations_q == (no_offset ? 1 : 0)) begin
            last_iteration_d = 1'b1;
            vrf_next_state = VRF_STORE_READ;
          // Send read request to memory
          end else begin
            num_iterations_d = num_iterations_q - 1;
            data_req_o = 1'b1;
            agu_get_rd_o = 1'b1;
            if (data_gnt_i) begin
              agu_incr_o = 1'b1;
              vrf_next_state = VRF_STORE_READ;
            end else begin
              vrf_next_state = VRF_STORE_WAITGNT;
            end
          end
        // we wait in this state
        end else begin
          vrf_next_state = VRF_STORE_WAITLSU;
        end
      end

      VRF_STORE_WAITGNT: begin
        data_req_o = 1'b1;
        agu_get_rd_o = 1'b1;
        if (data_gnt_i) begin
          agu_incr_o = 1'b1;
          vrf_next_state = VRF_STORE_READ;
        end else begin
          vrf_next_state = VRF_STORE_WAITGNT;
        end
      end

      // illegal state go back to idle
      default: begin
        vrf_next_state = VRF_IDLE;
      end
    endcase
  end

  ///////////////////////////
  // Delayed grant support //
  ///////////////////////////

  // Delayed read buffer
  assign rbuffer_d = rs1_d;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      curr_state_rdelay <= 1'b0;
      rbuffer_q <= '0;
    end else begin
      curr_state_rdelay <= next_state_rdelay;
      if (rbuffer_en) rbuffer_q <= rbuffer_d;
    end
  end
  always_comb begin
    rbuffer_en = 1'b0;
    case (curr_state_rdelay)
      1'b0: begin
        rdata_mux = 1'b0;
        if (read_delayed) begin
          rbuffer_en = 1'b1;
          next_state_rdelay = 1'b1;
        end else begin
          next_state_rdelay = 1'b0;
        end
      end
      1'b1: begin
        rdata_mux = 1'b1;
        if (read_delayed) begin
          next_state_rdelay = 1'b1;
        end else begin
          next_state_rdelay = 1'b0;
        end
      end
    endcase
  end

  // Delayed write buffer
  assign wbuffer_d = rd_q;
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      curr_state_wdelay <= 1'b0;
      wbuffer_q <= '0;
    end else begin
      curr_state_wdelay <= next_state_wdelay;
      if (wbuffer_en) wbuffer_q <= wbuffer_d;
    end
  end
  always_comb begin
    rd_buf_en = 1'b0;
    wbuffer_en = 1'b0;
    case (curr_state_wdelay)
      1'b0: begin
        wdata_mux = memory_op_i ? 2'b01 : 2'b00;
        if (write_delayed) begin
          if (!memory_op_i) rd_buf_en = 1'b1;
          else wbuffer_en = 1'b1;
          next_state_wdelay = 1'b1;
        end else begin
          next_state_wdelay = 1'b0;
        end
      end
      1'b1: begin
        wdata_mux = memory_op_i ? 2'b10 : 2'b01;
        if (write_delayed) begin
          next_state_wdelay = 1'b1;
        end else begin
          next_state_wdelay = 1'b0;
        end
      end
    endcase
  end

  ////////////////////////
  // Internal registers //
  ////////////////////////

  // Operands and result registers
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      rs1_q <= '0;
      rs2_q <= '0;
      rs3_q <= '0;
      rd_q  <= '0;
    end else begin
      if (rs1_en) rs1_q <= rs1_d;
      if (rs2_en) rs2_q <= rs2_d;
      if (rs3_en) rs3_q <= rs3_d;
      if (rd_en || rd_buf_en) rd_q <= rd_d;
    end
  end
  always_comb begin   // TODO: probably this condition is redundant and I should remove it
    rs1_d = rs1_en ? data_rdata_i : rs1_q;
    rs2_d = rs2_en ? data_rdata_i : rs2_q;
    rs3_d = rs3_en ? data_rdata_i : rs3_q;
    rd_d = wdata_i;
  end

  /////////////
  // Outputs //
  /////////////

  assign rdata_a_o = rdata_mux ? rbuffer_q : rs1_q;
  assign rdata_b_o = rs2_q;
  assign rdata_c_o = rs3_q;
  // mux for the write data
  always_comb begin
    case (wdata_mux)
      2'b00: data_wdata_o = wdata_i;
      2'b01: data_wdata_o = rd_q;
      2'b10: data_wdata_o = wbuffer_q;
      default: data_wdata_o = '0;
    endcase
  end

endmodule
